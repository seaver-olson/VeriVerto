module alu(input wire[31:0] A, input wire[31:0] B, input wire[7:0]);
    
endmodule