module IF_ID(
    input wire [31:0] instruction,
    input wire [31:0] pc,
    input wire writeFlag,
    output wire [31:0] instruction
);

endmodule