module EX_MEM(

);

endmodule