module equalityTestUnit();

endmodule