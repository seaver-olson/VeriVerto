module pcUnit(
    input wire clk,
    input wire rst,
    inp
);
    wire [31:0] pcIncr;
    
endmodule