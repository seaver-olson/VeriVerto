module hazardDetectionUnit(
    
);

endmodule