module regfile(input clk);
    //sync clock to io exec
    always @(posedge clk) begin
        
    end
endmodule