module ID_EX(

);

endmodule