module forwardingUnit(
    input wire [31:0] EX_MEM_writeReg
    input wire [31:0] MEM_WB_writeReg,
    output wire [1:0] ForwardA,
    output wire [1:0] FordwardB
);

endmodule