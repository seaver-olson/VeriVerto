module MEM_WB(

);

endmodule